import CacheTypes::*;
import Vector::*;
import MemTypes::*;
import Types::*;
import ProcTypes::*;
import Fifo::*;
import Ehr::*;

// TODO: implement I cache for Ex 1

module mkICache(WideMem mem, ICache ifc);

endmodule

